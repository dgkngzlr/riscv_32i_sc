----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:44:09 06/10/2022 
-- Design Name: 
-- Module Name:    div - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity div is
port(
	i_en: in std_logic;
	i_a : in std_logic_vector(31 downto 0);
	i_b : in std_logic_vector(31 downto 0);
	o_r : out std_logic_vector(31 downto 0)
);
end div;

architecture Behavioral of div is

begin

process(i_a, i_b, i_en)
begin
	if i_en = '1' and i_b /= x"00000000" then
		o_r <= std_logic_vector(unsigned(i_a) / unsigned(i_b));
	else
		o_r <= (others => '0');
	end if;
end process;

end Behavioral;

